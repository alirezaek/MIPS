library verilog;
use verilog.vl_types.all;
entity Mux32bit_tb is
end Mux32bit_tb;
