library verilog;
use verilog.vl_types.all;
entity CPU_Core is
    port(
        clk             : in     vl_logic
    );
end CPU_Core;
