/*
  MIPS SINGLE CYCLE CPU IMPLEMENTED BY :   
  ARDESHIR  ALIREZA 
  92213118  92213034
*/
module PC (
  input in,
  output out
  );
  
  assign out = in;
  
endmodule
