library verilog;
use verilog.vl_types.all;
entity PC is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end PC;
