library verilog;
use verilog.vl_types.all;
entity Test is
    port(
        in1             : in     vl_logic_vector(31 downto 0);
        \out\           : out    vl_logic_vector(34 downto 0)
    );
end Test;
