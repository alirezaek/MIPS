library verilog;
use verilog.vl_types.all;
entity Test_Bench2 is
end Test_Bench2;
